module sample (
	a,
	b,
	c, d, e
);
input [7:0] a, b, c;
output d, e;

reg	hoge, _dff123;


endmodule
