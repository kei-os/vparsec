module sample;endmodule
