module sample(a);

input a;

reg b[1:0], c;
reg [1:0] d, e[3:0], f;

endmodule
