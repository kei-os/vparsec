module sample (
	a,
	b,
	c
);
input [:] a, b, c;


endmodule
