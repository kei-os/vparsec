module sample (
	a,
	b,
	c
);

endmodule
